LIBRARY ieee;